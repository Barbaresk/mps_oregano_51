
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;
LIBRARY UNISIM;
USE UNISIM.Vcomponents.ALL;
ENTITY top_mps_top_mps_sch_tb IS
END top_mps_top_mps_sch_tb;
ARCHITECTURE behavioral OF top_mps_top_mps_sch_tb IS 

   COMPONENT top_mps
   PORT( RESET	:	IN	STD_LOGIC; 
          RAMX_ACCESS_EN	:	IN	STD_LOGIC; 
          RAMX_DATA_VALID	:	IN	STD_LOGIC; 
          INT0_I	:	IN	STD_LOGIC_VECTOR (0 DOWNTO 0); 
          INT1_I	:	IN	STD_LOGIC_VECTOR (0 DOWNTO 0); 
          ALL_T0_I	:	IN	STD_LOGIC_VECTOR (0 DOWNTO 0); 
          ALL_T1_I	:	IN	STD_LOGIC_VECTOR (0 DOWNTO 0); 
          ALL_RXD_I	:	IN	STD_LOGIC_VECTOR (0 DOWNTO 0); 
          P0_I	:	IN	STD_LOGIC_VECTOR (7 DOWNTO 0); 
          P1_I	:	IN	STD_LOGIC_VECTOR (7 DOWNTO 0); 
          P2_I	:	IN	STD_LOGIC_VECTOR (7 DOWNTO 0); 
          P3_I	:	IN	STD_LOGIC_VECTOR (7 DOWNTO 0); 
          RAMX_RD	:	OUT	STD_LOGIC; 
          P0_O	:	OUT	STD_LOGIC_VECTOR (7 DOWNTO 0); 
          P1_O	:	OUT	STD_LOGIC_VECTOR (7 DOWNTO 0); 
          P2_O	:	OUT	STD_LOGIC_VECTOR (7 DOWNTO 0); 
          P3_O	:	OUT	STD_LOGIC_VECTOR (7 DOWNTO 0); 
          ALL_RXD_O	:	OUT	STD_LOGIC_VECTOR (0 DOWNTO 0); 
          ALL_TXD_O	:	OUT	STD_LOGIC_VECTOR (0 DOWNTO 0); 
          ALL_RXDWR_O	:	OUT	STD_LOGIC_VECTOR (0 DOWNTO 0); 
          CLK	:	IN	STD_LOGIC; 
          LOAD	:	IN	STD_LOGIC; 
          UD	:	IN	STD_LOGIC; 
          COUNT	:	IN	STD_LOGIC_VECTOR (7 DOWNTO 0));
   END COMPONENT;

   SIGNAL RESET	:	STD_LOGIC := '0';
   SIGNAL RAMX_ACCESS_EN	:	STD_LOGIC := '0';
   SIGNAL RAMX_DATA_VALID	:	STD_LOGIC := '0';
   SIGNAL INT0_I	:	STD_LOGIC_VECTOR (0 DOWNTO 0) := "0";
   SIGNAL INT1_I	:	STD_LOGIC_VECTOR (0 DOWNTO 0) := "0";
   SIGNAL ALL_T0_I	:	STD_LOGIC_VECTOR (0 DOWNTO 0) := "0";
   SIGNAL ALL_T1_I	:	STD_LOGIC_VECTOR (0 DOWNTO 0) := "0";
   SIGNAL ALL_RXD_I	:	STD_LOGIC_VECTOR (0 DOWNTO 0) := "0";
   SIGNAL P0_I	:	STD_LOGIC_VECTOR (7 DOWNTO 0) := (others => '0');
   SIGNAL P1_I	:	STD_LOGIC_VECTOR (7 DOWNTO 0) := (others => '0');
   SIGNAL P2_I	:	STD_LOGIC_VECTOR (7 DOWNTO 0) := (others => '0');
   SIGNAL P3_I	:	STD_LOGIC_VECTOR (7 DOWNTO 0) := (others => '0');
   SIGNAL RAMX_RD	:	STD_LOGIC;
   SIGNAL P0_O	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
   SIGNAL P1_O	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
   SIGNAL P2_O	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
   SIGNAL P3_O	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
   SIGNAL ALL_RXD_O	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
   SIGNAL ALL_TXD_O	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
   SIGNAL ALL_RXDWR_O	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
   SIGNAL CLK	:	STD_LOGIC := '0';
   SIGNAL LOAD	:	STD_LOGIC := '0';
   SIGNAL UD	:	STD_LOGIC := '0';
   SIGNAL COUNT	:	STD_LOGIC_VECTOR (7 DOWNTO 0) := (others => '0');

	constant CLK_T : time := 10 ns;
BEGIN

   UUT: top_mps PORT MAP(
		RESET => RESET, 
		RAMX_ACCESS_EN => RAMX_ACCESS_EN, 
		RAMX_DATA_VALID => RAMX_DATA_VALID, 
		INT0_I => INT0_I, 
		INT1_I => INT1_I, 
		ALL_T0_I => ALL_T0_I, 
		ALL_T1_I => ALL_T1_I, 
		ALL_RXD_I => ALL_RXD_I, 
		P0_I => P0_I, 
		P1_I => P1_I, 
		P2_I => P2_I, 
		P3_I => P3_I, 
		RAMX_RD => RAMX_RD, 
		P0_O => P0_O, 
		P1_O => P1_O, 
		P2_O => P2_O, 
		P3_O => P3_O, 
		ALL_RXD_O => ALL_RXD_O, 
		ALL_TXD_O => ALL_TXD_O, 
		ALL_RXDWR_O => ALL_RXDWR_O, 
		CLK => CLK, 
		LOAD => LOAD, 
		UD => UD, 
		COUNT => COUNT
   );
	
	CLK <= not CLK after CLK_T / 2;
	process begin
		RESET <= '1';
		wait for 40 * CLK_T;
		RESET <= '0';
		RAMX_ACCESS_EN <= '1';
		wait for 100 * CLK_T;
	
	end process;

END;